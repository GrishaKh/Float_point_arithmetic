module round (exp, mantis, sign, operator, loss, mantis_out, exp_out);

input sign;
input [7:0] exp;
input [27:0] mantis;
input loss;
input operator;
output [7:0] exp_out;
output [22:0] mantis_out;

wire [23:0] mantis_tmp;
wire carry;
wire [3:0] r_bits = mantis[3:0];
wire [27:0] mantis_shifted;

assign exp_out = exp;
//assign mantis_out = mantis_shifted[26:4];
assign mantis_out = |exp ? mantis_tmp[22:0] : mantis_tmp[23:1];

//assign {carry, mantis_tmp} = mantis[3:0] > 4'b1000 ? 
//				mantis[26:4] + mantis[3] : mantis[26:4];

assign {carry, mantis_tmp} = (r_bits > 4'b1000 || (r_bits == 4'b1000 && mantis[4] | loss)) ?
			mantis[27:4] + mantis[3] : mantis[27:4];

/*always @(*) begin
    if (operator) begin
        if (r_bits < 4'b1000) 
    end
end*/

/*shifter #(.DIRECTION(1)) __shifter (
    .exp (exp),
    .exp_target_or_diff ({{7{1'b0}}, carry}),
    .mantis (mantis_tmp),
    .exp_out (exp_out),
    .mantis_out (mantis_shifted)
);*/

endmodule // round
