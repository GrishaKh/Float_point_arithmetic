module standardizer (
    exp_in, mantis_in,
    exp_out, mantis_out
);

input [7:0] exp_in;
input [27:0] mantis_in;
output [7:0] exp_out
output [22:0] mantis_out;



endmodule // standardizer