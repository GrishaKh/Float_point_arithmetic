module preadder (
    number_A, number_B,
    sign, exp,
    mantis_great, mantis_small
);

endmodule // preadder